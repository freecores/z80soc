library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
        port(
                Clk : in std_logic;
                A   : in std_logic_vector(13 downto 0);
                D   : out std_logic_vector(7 downto 0)
        );
end rom;

architecture rtl of rom is
begin

process (Clk)
begin
 if Clk'event and Clk = '1' then
        case A is
             when "00000000000000" => D <= x"ED";
             when "00000000000001" => D <= x"7B";
             when "00000000000010" => D <= x"DE";
             when "00000000000011" => D <= x"7F";
             when "00000000000100" => D <= x"3A";
             when "00000000000101" => D <= x"DD";
             when "00000000000110" => D <= x"7F";
             when "00000000000111" => D <= x"B7";
             when "00000000001000" => D <= x"28";
             when "00000000001001" => D <= x"03";
             when "00000000001010" => D <= x"CD";
             when "00000000001011" => D <= x"96";
             when "00000000001100" => D <= x"01";
             when "00000000001101" => D <= x"CD";
             when "00000000001110" => D <= x"F4";
             when "00000000001111" => D <= x"00";
             when "00000000010000" => D <= x"11";
             when "00000000010001" => D <= x"34";
             when "00000000010010" => D <= x"40";
             when "00000000010011" => D <= x"21";
             when "00000000010100" => D <= x"12";
             when "00000000010101" => D <= x"02";
             when "00000000010110" => D <= x"CD";
             when "00000000010111" => D <= x"07";
             when "00000000011000" => D <= x"01";
             when "00000000011001" => D <= x"11";
             when "00000000011010" => D <= x"5C";
             when "00000000011011" => D <= x"40";
             when "00000000011100" => D <= x"21";
             when "00000000011101" => D <= x"25";
             when "00000000011110" => D <= x"02";
             when "00000000011111" => D <= x"CD";
             when "00000000100000" => D <= x"07";
             when "00000000100001" => D <= x"01";
             when "00000000100010" => D <= x"CD";
             when "00000000100011" => D <= x"12";
             when "00000000100100" => D <= x"01";
             when "00000000100101" => D <= x"11";
             when "00000000100110" => D <= x"46";
             when "00000000100111" => D <= x"41";
             when "00000000101000" => D <= x"21";
             when "00000000101001" => D <= x"38";
             when "00000000101010" => D <= x"02";
             when "00000000101011" => D <= x"CD";
             when "00000000101100" => D <= x"07";
             when "00000000101101" => D <= x"01";
             when "00000000101110" => D <= x"11";
             when "00000000101111" => D <= x"96";
             when "00000000110000" => D <= x"41";
             when "00000000110001" => D <= x"21";
             when "00000000110010" => D <= x"54";
             when "00000000110011" => D <= x"02";
             when "00000000110100" => D <= x"CD";
             when "00000000110101" => D <= x"07";
             when "00000000110110" => D <= x"01";
             when "00000000110111" => D <= x"11";
             when "00000000111000" => D <= x"E6";
             when "00000000111001" => D <= x"41";
             when "00000000111010" => D <= x"21";
             when "00000000111011" => D <= x"71";
             when "00000000111100" => D <= x"02";
             when "00000000111101" => D <= x"CD";
             when "00000000111110" => D <= x"07";
             when "00000000111111" => D <= x"01";
             when "00000001000000" => D <= x"11";
             when "00000001000001" => D <= x"36";
             when "00000001000010" => D <= x"42";
             when "00000001000011" => D <= x"21";
             when "00000001000100" => D <= x"8E";
             when "00000001000101" => D <= x"02";
             when "00000001000110" => D <= x"CD";
             when "00000001000111" => D <= x"07";
             when "00000001001000" => D <= x"01";
             when "00000001001001" => D <= x"11";
             when "00000001001010" => D <= x"5E";
             when "00000001001011" => D <= x"42";
             when "00000001001100" => D <= x"21";
             when "00000001001101" => D <= x"A2";
             when "00000001001110" => D <= x"02";
             when "00000001001111" => D <= x"CD";
             when "00000001010000" => D <= x"07";
             when "00000001010001" => D <= x"01";
             when "00000001010010" => D <= x"21";
             when "00000001010011" => D <= x"45";
             when "00000001010100" => D <= x"03";
             when "00000001010101" => D <= x"3A";
             when "00000001010110" => D <= x"DD";
             when "00000001010111" => D <= x"7F";
             when "00000001011000" => D <= x"B7";
             when "00000001011001" => D <= x"28";
             when "00000001011010" => D <= x"03";
             when "00000001011011" => D <= x"21";
             when "00000001011100" => D <= x"51";
             when "00000001011101" => D <= x"03";
             when "00000001011110" => D <= x"11";
             when "00000001011111" => D <= x"87";
             when "00000001100000" => D <= x"40";
             when "00000001100001" => D <= x"CD";
             when "00000001100010" => D <= x"07";
             when "00000001100011" => D <= x"01";
             when "00000001100100" => D <= x"11";
             when "00000001100101" => D <= x"D6";
             when "00000001100110" => D <= x"42";
             when "00000001100111" => D <= x"01";
             when "00000001101000" => D <= x"1E";
             when "00000001101001" => D <= x"00";
             when "00000001101010" => D <= x"C5";
             when "00000001101011" => D <= x"D5";
             when "00000001101100" => D <= x"CD";
             when "00000001101101" => D <= x"DF";
             when "00000001101110" => D <= x"00";
             when "00000001101111" => D <= x"CD";
             when "00000001110000" => D <= x"3C";
             when "00000001110001" => D <= x"01";
             when "00000001110010" => D <= x"3A";
             when "00000001110011" => D <= x"DD";
             when "00000001110100" => D <= x"7F";
             when "00000001110101" => D <= x"B7";
             when "00000001110110" => D <= x"28";
             when "00000001110111" => D <= x"03";
             when "00000001111000" => D <= x"CD";
             when "00000001111001" => D <= x"6F";
             when "00000001111010" => D <= x"01";
             when "00000001111011" => D <= x"CD";
             when "00000001111100" => D <= x"0F";
             when "00000001111101" => D <= x"01";
             when "00000001111110" => D <= x"D1";
             when "00000001111111" => D <= x"C1";
             when "00000010000000" => D <= x"B7";
             when "00000010000001" => D <= x"28";
             when "00000010000010" => D <= x"E7";
             when "00000010000011" => D <= x"FE";
             when "00000010000100" => D <= x"41";
             when "00000010000101" => D <= x"28";
             when "00000010000110" => D <= x"15";
             when "00000010000111" => D <= x"D3";
             when "00000010001000" => D <= x"01";
             when "00000010001001" => D <= x"6F";
             when "00000010001010" => D <= x"3A";
             when "00000010001011" => D <= x"DD";
             when "00000010001100" => D <= x"7F";
             when "00000010001101" => D <= x"B7";
             when "00000010001110" => D <= x"20";
             when "00000010001111" => D <= x"03";
             when "00000010010000" => D <= x"7D";
             when "00000010010001" => D <= x"D3";
             when "00000010010010" => D <= x"11";
             when "00000010010011" => D <= x"12";
             when "00000010010100" => D <= x"13";
             when "00000010010101" => D <= x"0B";
             when "00000010010110" => D <= x"78";
             when "00000010010111" => D <= x"B1";
             when "00000010011000" => D <= x"28";
             when "00000010011001" => D <= x"CA";
             when "00000010011010" => D <= x"18";
             when "00000010011011" => D <= x"CE";
             when "00000010011100" => D <= x"21";
             when "00000010011101" => D <= x"00";
             when "00000010011110" => D <= x"80";
             when "00000010011111" => D <= x"3E";
             when "00000010100000" => D <= x"00";
             when "00000010100001" => D <= x"77";
             when "00000010100010" => D <= x"23";
             when "00000010100011" => D <= x"3C";
             when "00000010100100" => D <= x"20";
             when "00000010100101" => D <= x"FB";
             when "00000010100110" => D <= x"CD";
             when "00000010100111" => D <= x"CA";
             when "00000010101000" => D <= x"00";
             when "00000010101001" => D <= x"21";
             when "00000010101010" => D <= x"00";
             when "00000010101011" => D <= x"80";
             when "00000010101100" => D <= x"3A";
             when "00000010101101" => D <= x"DD";
             when "00000010101110" => D <= x"7F";
             when "00000010101111" => D <= x"B7";
             when "00000010110000" => D <= x"20";
             when "00000010110001" => D <= x"06";
             when "00000010110010" => D <= x"7C";
             when "00000010110011" => D <= x"D3";
             when "00000010110100" => D <= x"11";
             when "00000010110101" => D <= x"7D";
             when "00000010110110" => D <= x"D3";
             when "00000010110111" => D <= x"10";
             when "00000010111000" => D <= x"7E";
             when "00000010111001" => D <= x"D3";
             when "00000010111010" => D <= x"01";
             when "00000010111011" => D <= x"CD";
             when "00000010111100" => D <= x"DF";
             when "00000010111101" => D <= x"00";
             when "00000010111110" => D <= x"23";
             when "00000010111111" => D <= x"7E";
             when "00000011000000" => D <= x"FE";
             when "00000011000001" => D <= x"FF";
             when "00000011000010" => D <= x"20";
             when "00000011000011" => D <= x"F4";
             when "00000011000100" => D <= x"CD";
             when "00000011000101" => D <= x"CA";
             when "00000011000110" => D <= x"00";
             when "00000011000111" => D <= x"C3";
             when "00000011001000" => D <= x"04";
             when "00000011001001" => D <= x"00";
             when "00000011001010" => D <= x"CD";
             when "00000011001011" => D <= x"DF";
             when "00000011001100" => D <= x"00";
             when "00000011001101" => D <= x"DB";
             when "00000011001110" => D <= x"30";
             when "00000011001111" => D <= x"FE";
             when "00000011010000" => D <= x"01";
             when "00000011010001" => D <= x"20";
             when "00000011010010" => D <= x"F7";
             when "00000011010011" => D <= x"C9";
             when "00000011010100" => D <= x"DB";
             when "00000011010101" => D <= x"20";
             when "00000011010110" => D <= x"B7";
             when "00000011010111" => D <= x"20";
             when "00000011011000" => D <= x"02";
             when "00000011011001" => D <= x"3E";
             when "00000011011010" => D <= x"01";
             when "00000011011011" => D <= x"3D";
             when "00000011011100" => D <= x"20";
             when "00000011011101" => D <= x"FD";
             when "00000011011110" => D <= x"C9";
             when "00000011011111" => D <= x"DB";
             when "00000011100000" => D <= x"20";
             when "00000011100001" => D <= x"B7";
             when "00000011100010" => D <= x"20";
             when "00000011100011" => D <= x"02";
             when "00000011100100" => D <= x"3E";
             when "00000011100101" => D <= x"01";
             when "00000011100110" => D <= x"F5";
             when "00000011100111" => D <= x"01";
             when "00000011101000" => D <= x"88";
             when "00000011101001" => D <= x"13";
             when "00000011101010" => D <= x"0B";
             when "00000011101011" => D <= x"78";
             when "00000011101100" => D <= x"B1";
             when "00000011101101" => D <= x"20";
             when "00000011101110" => D <= x"FB";
             when "00000011101111" => D <= x"F1";
             when "00000011110000" => D <= x"3D";
             when "00000011110001" => D <= x"20";
             when "00000011110010" => D <= x"F3";
             when "00000011110011" => D <= x"C9";
             when "00000011110100" => D <= x"3E";
             when "00000011110101" => D <= x"00";
             when "00000011110110" => D <= x"D3";
             when "00000011110111" => D <= x"91";
             when "00000011111000" => D <= x"D3";
             when "00000011111001" => D <= x"92";
             when "00000011111010" => D <= x"01";
             when "00000011111011" => D <= x"B0";
             when "00000011111100" => D <= x"04";
             when "00000011111101" => D <= x"3E";
             when "00000011111110" => D <= x"20";
             when "00000011111111" => D <= x"D3";
             when "00000100000000" => D <= x"90";
             when "00000100000001" => D <= x"0B";
             when "00000100000010" => D <= x"78";
             when "00000100000011" => D <= x"B1";
             when "00000100000100" => D <= x"20";
             when "00000100000101" => D <= x"F7";
             when "00000100000110" => D <= x"C9";
             when "00000100000111" => D <= x"7E";
             when "00000100001000" => D <= x"B7";
             when "00000100001001" => D <= x"C8";
             when "00000100001010" => D <= x"12";
             when "00000100001011" => D <= x"23";
             when "00000100001100" => D <= x"13";
             when "00000100001101" => D <= x"18";
             when "00000100001110" => D <= x"F8";
             when "00000100001111" => D <= x"DB";
             when "00000100010000" => D <= x"80";
             when "00000100010001" => D <= x"C9";
             when "00000100010010" => D <= x"21";
             when "00000100010011" => D <= x"C1";
             when "00000100010100" => D <= x"02";
             when "00000100010101" => D <= x"11";
             when "00000100010110" => D <= x"F5";
             when "00000100010111" => D <= x"40";
             when "00000100011000" => D <= x"CD";
             when "00000100011001" => D <= x"07";
             when "00000100011010" => D <= x"01";
             when "00000100011011" => D <= x"11";
             when "00000100011100" => D <= x"1D";
             when "00000100011101" => D <= x"41";
             when "00000100011110" => D <= x"3E";
             when "00000100011111" => D <= x"0A";
             when "00000100100000" => D <= x"21";
             when "00000100100001" => D <= x"03";
             when "00000100100010" => D <= x"03";
             when "00000100100011" => D <= x"E5";
             when "00000100100100" => D <= x"F5";
             when "00000100100101" => D <= x"D5";
             when "00000100100110" => D <= x"CD";
             when "00000100100111" => D <= x"07";
             when "00000100101000" => D <= x"01";
             when "00000100101001" => D <= x"D1";
             when "00000100101010" => D <= x"F1";
             when "00000100101011" => D <= x"21";
             when "00000100101100" => D <= x"28";
             when "00000100101101" => D <= x"00";
             when "00000100101110" => D <= x"19";
             when "00000100101111" => D <= x"54";
             when "00000100110000" => D <= x"5D";
             when "00000100110001" => D <= x"E1";
             when "00000100110010" => D <= x"3D";
             when "00000100110011" => D <= x"20";
             when "00000100110100" => D <= x"EB";
             when "00000100110101" => D <= x"21";
             when "00000100110110" => D <= x"E2";
             when "00000100110111" => D <= x"02";
             when "00000100111000" => D <= x"CD";
             when "00000100111001" => D <= x"07";
             when "00000100111010" => D <= x"01";
             when "00000100111011" => D <= x"C9";
             when "00000100111100" => D <= x"21";
             when "00000100111101" => D <= x"1E";
             when "00000100111110" => D <= x"41";
             when "00000100111111" => D <= x"11";
             when "00000101000000" => D <= x"00";
             when "00000101000001" => D <= x"90";
             when "00000101000010" => D <= x"01";
             when "00000101000011" => D <= x"1E";
             when "00000101000100" => D <= x"00";
             when "00000101000101" => D <= x"ED";
             when "00000101000110" => D <= x"B0";
             when "00000101000111" => D <= x"21";
             when "00000101001000" => D <= x"46";
             when "00000101001001" => D <= x"41";
             when "00000101001010" => D <= x"11";
             when "00000101001011" => D <= x"1E";
             when "00000101001100" => D <= x"41";
             when "00000101001101" => D <= x"06";
             when "00000101001110" => D <= x"09";
             when "00000101001111" => D <= x"C5";
             when "00000101010000" => D <= x"E5";
             when "00000101010001" => D <= x"D5";
             when "00000101010010" => D <= x"01";
             when "00000101010011" => D <= x"1E";
             when "00000101010100" => D <= x"00";
             when "00000101010101" => D <= x"ED";
             when "00000101010110" => D <= x"B0";
             when "00000101010111" => D <= x"D1";
             when "00000101011000" => D <= x"21";
             when "00000101011001" => D <= x"28";
             when "00000101011010" => D <= x"00";
             when "00000101011011" => D <= x"19";
             when "00000101011100" => D <= x"54";
             when "00000101011101" => D <= x"5D";
             when "00000101011110" => D <= x"E1";
             when "00000101011111" => D <= x"01";
             when "00000101100000" => D <= x"28";
             when "00000101100001" => D <= x"00";
             when "00000101100010" => D <= x"09";
             when "00000101100011" => D <= x"C1";
             when "00000101100100" => D <= x"10";
             when "00000101100101" => D <= x"E9";
             when "00000101100110" => D <= x"21";
             when "00000101100111" => D <= x"00";
             when "00000101101000" => D <= x"90";
             when "00000101101001" => D <= x"01";
             when "00000101101010" => D <= x"1E";
             when "00000101101011" => D <= x"00";
             when "00000101101100" => D <= x"ED";
             when "00000101101101" => D <= x"B0";
             when "00000101101110" => D <= x"C9";
             when "00000101101111" => D <= x"C5";
             when "00000101110000" => D <= x"D5";
             when "00000101110001" => D <= x"CD";
             when "00000101110010" => D <= x"AD";
             when "00000101110011" => D <= x"01";
             when "00000101110100" => D <= x"FE";
             when "00000101110101" => D <= x"01";
             when "00000101110110" => D <= x"20";
             when "00000101110111" => D <= x"07";
             when "00000101111000" => D <= x"CD";
             when "00000101111001" => D <= x"EE";
             when "00000101111010" => D <= x"01";
             when "00000101111011" => D <= x"3E";
             when "00000101111100" => D <= x"01";
             when "00000101111101" => D <= x"18";
             when "00000101111110" => D <= x"09";
             when "00000101111111" => D <= x"FE";
             when "00000110000000" => D <= x"02";
             when "00000110000001" => D <= x"20";
             when "00000110000010" => D <= x"10";
             when "00000110000011" => D <= x"CD";
             when "00000110000100" => D <= x"CA";
             when "00000110000101" => D <= x"01";
             when "00000110000110" => D <= x"3E";
             when "00000110000111" => D <= x"80";
             when "00000110001000" => D <= x"D3";
             when "00000110001001" => D <= x"01";
             when "00000110001010" => D <= x"11";
             when "00000110001011" => D <= x"E0";
             when "00000110001100" => D <= x"7F";
             when "00000110001101" => D <= x"21";
             when "00000110001110" => D <= x"00";
             when "00000110001111" => D <= x"91";
             when "00000110010000" => D <= x"CD";
             when "00000110010001" => D <= x"07";
             when "00000110010010" => D <= x"01";
             when "00000110010011" => D <= x"D1";
             when "00000110010100" => D <= x"C1";
             when "00000110010101" => D <= x"C9";
             when "00000110010110" => D <= x"11";
             when "00000110010111" => D <= x"00";
             when "00000110011000" => D <= x"91";
             when "00000110011001" => D <= x"21";
             when "00000110011010" => D <= x"24";
             when "00000110011011" => D <= x"03";
             when "00000110011100" => D <= x"01";
             when "00000110011101" => D <= x"21";
             when "00000110011110" => D <= x"00";
             when "00000110011111" => D <= x"ED";
             when "00000110100000" => D <= x"B0";
             when "00000110100001" => D <= x"11";
             when "00000110100010" => D <= x"E0";
             when "00000110100011" => D <= x"7F";
             when "00000110100100" => D <= x"21";
             when "00000110100101" => D <= x"00";
             when "00000110100110" => D <= x"91";
             when "00000110100111" => D <= x"01";
             when "00000110101000" => D <= x"20";
             when "00000110101001" => D <= x"00";
             when "00000110101010" => D <= x"ED";
             when "00000110101011" => D <= x"B0";
             when "00000110101100" => D <= x"C9";
             when "00000110101101" => D <= x"CD";
             when "00000110101110" => D <= x"BE";
             when "00000110101111" => D <= x"01";
             when "00000110110000" => D <= x"3E";
             when "00000110110001" => D <= x"00";
             when "00000110110010" => D <= x"C0";
             when "00000110110011" => D <= x"DB";
             when "00000110110100" => D <= x"70";
             when "00000110110101" => D <= x"C9";
             when "00000110110110" => D <= x"3A";
             when "00000110110111" => D <= x"00";
             when "00000110111000" => D <= x"90";
             when "00000110111001" => D <= x"3D";
             when "00000110111010" => D <= x"32";
             when "00000110111011" => D <= x"00";
             when "00000110111100" => D <= x"90";
             when "00000110111101" => D <= x"C9";
             when "00000110111110" => D <= x"3A";
             when "00000110111111" => D <= x"01";
             when "00000111000000" => D <= x"90";
             when "00000111000001" => D <= x"3D";
             when "00000111000010" => D <= x"20";
             when "00000111000011" => D <= x"02";
             when "00000111000100" => D <= x"3E";
             when "00000111000101" => D <= x"10";
             when "00000111000110" => D <= x"32";
             when "00000111000111" => D <= x"01";
             when "00000111001000" => D <= x"90";
             when "00000111001001" => D <= x"C9";
             when "00000111001010" => D <= x"3A";
             when "00000111001011" => D <= x"00";
             when "00000111001100" => D <= x"91";
             when "00000111001101" => D <= x"32";
             when "00000111001110" => D <= x"02";
             when "00000111001111" => D <= x"90";
             when "00000111010000" => D <= x"3A";
             when "00000111010001" => D <= x"10";
             when "00000111010010" => D <= x"91";
             when "00000111010011" => D <= x"32";
             when "00000111010100" => D <= x"03";
             when "00000111010101" => D <= x"90";
             when "00000111010110" => D <= x"21";
             when "00000111010111" => D <= x"01";
             when "00000111011000" => D <= x"91";
             when "00000111011001" => D <= x"11";
             when "00000111011010" => D <= x"00";
             when "00000111011011" => D <= x"91";
             when "00000111011100" => D <= x"01";
             when "00000111011101" => D <= x"1F";
             when "00000111011110" => D <= x"00";
             when "00000111011111" => D <= x"ED";
             when "00000111100000" => D <= x"B0";
             when "00000111100001" => D <= x"3A";
             when "00000111100010" => D <= x"02";
             when "00000111100011" => D <= x"90";
             when "00000111100100" => D <= x"32";
             when "00000111100101" => D <= x"0F";
             when "00000111100110" => D <= x"91";
             when "00000111100111" => D <= x"3A";
             when "00000111101000" => D <= x"03";
             when "00000111101001" => D <= x"90";
             when "00000111101010" => D <= x"32";
             when "00000111101011" => D <= x"1F";
             when "00000111101100" => D <= x"91";
             when "00000111101101" => D <= x"C9";
             when "00000111101110" => D <= x"3A";
             when "00000111101111" => D <= x"0F";
             when "00000111110000" => D <= x"91";
             when "00000111110001" => D <= x"32";
             when "00000111110010" => D <= x"02";
             when "00000111110011" => D <= x"90";
             when "00000111110100" => D <= x"3A";
             when "00000111110101" => D <= x"1F";
             when "00000111110110" => D <= x"91";
             when "00000111110111" => D <= x"32";
             when "00000111111000" => D <= x"03";
             when "00000111111001" => D <= x"90";
             when "00000111111010" => D <= x"21";
             when "00000111111011" => D <= x"1E";
             when "00000111111100" => D <= x"91";
             when "00000111111101" => D <= x"11";
             when "00000111111110" => D <= x"1F";
             when "00000111111111" => D <= x"91";
             when "00001000000000" => D <= x"01";
             when "00001000000001" => D <= x"1F";
             when "00001000000010" => D <= x"00";
             when "00001000000011" => D <= x"ED";
             when "00001000000100" => D <= x"B8";
             when "00001000000101" => D <= x"3A";
             when "00001000000110" => D <= x"02";
             when "00001000000111" => D <= x"90";
             when "00001000001000" => D <= x"32";
             when "00001000001001" => D <= x"00";
             when "00001000001010" => D <= x"91";
             when "00001000001011" => D <= x"3A";
             when "00001000001100" => D <= x"03";
             when "00001000001101" => D <= x"90";
             when "00001000001110" => D <= x"32";
             when "00001000001111" => D <= x"10";
             when "00001000010000" => D <= x"91";
             when "00001000010001" => D <= x"C9";
             when "00001000010010" => D <= x"5A";
             when "00001000010011" => D <= x"38";
             when "00001000010100" => D <= x"30";
             when "00001000010101" => D <= x"20";
             when "00001000010110" => D <= x"53";
             when "00001000010111" => D <= x"59";
             when "00001000011000" => D <= x"53";
             when "00001000011001" => D <= x"54";
             when "00001000011010" => D <= x"45";
             when "00001000011011" => D <= x"4D";
             when "00001000011100" => D <= x"20";
             when "00001000011101" => D <= x"4F";
             when "00001000011110" => D <= x"4E";
             when "00001000011111" => D <= x"20";
             when "00001000100000" => D <= x"43";
             when "00001000100001" => D <= x"48";
             when "00001000100010" => D <= x"49";
             when "00001000100011" => D <= x"50";
             when "00001000100100" => D <= x"00";
             when "00001000100101" => D <= x"52";
             when "00001000100110" => D <= x"4F";
             when "00001000100111" => D <= x"4E";
             when "00001000101000" => D <= x"49";
             when "00001000101001" => D <= x"56";
             when "00001000101010" => D <= x"4F";
             when "00001000101011" => D <= x"4E";
             when "00001000101100" => D <= x"20";
             when "00001000101101" => D <= x"43";
             when "00001000101110" => D <= x"4F";
             when "00001000101111" => D <= x"53";
             when "00001000110000" => D <= x"54";
             when "00001000110001" => D <= x"41";
             when "00001000110010" => D <= x"20";
             when "00001000110011" => D <= x"32";
             when "00001000110100" => D <= x"30";
             when "00001000110101" => D <= x"30";
             when "00001000110110" => D <= x"38";
             when "00001000110111" => D <= x"00";
             when "00001000111000" => D <= x"20";
             when "00001000111001" => D <= x"20";
             when "00001000111010" => D <= x"7C";
             when "00001000111011" => D <= x"21";
             when "00001000111100" => D <= x"23";
             when "00001000111101" => D <= x"24";
             when "00001000111110" => D <= x"25";
             when "00001000111111" => D <= x"26";
             when "00001001000000" => D <= x"2F";
             when "00001001000001" => D <= x"28";
             when "00001001000010" => D <= x"29";
             when "00001001000011" => D <= x"3D";
             when "00001001000100" => D <= x"3F";
             when "00001001000101" => D <= x"2A";
             when "00001001000110" => D <= x"60";
             when "00001001000111" => D <= x"2B";
             when "00001001001000" => D <= x"B4";
             when "00001001001001" => D <= x"E7";
             when "00001001001010" => D <= x"7E";
             when "00001001001011" => D <= x"5E";
             when "00001001001100" => D <= x"2C";
             when "00001001001101" => D <= x"2E";
             when "00001001001110" => D <= x"3B";
             when "00001001001111" => D <= x"3A";
             when "00001001010000" => D <= x"5C";
             when "00001001010001" => D <= x"3C";
             when "00001001010010" => D <= x"3E";
             when "00001001010011" => D <= x"00";
             when "00001001010100" => D <= x"20";
             when "00001001010101" => D <= x"20";
             when "00001001010110" => D <= x"41";
             when "00001001010111" => D <= x"42";
             when "00001001011000" => D <= x"43";
             when "00001001011001" => D <= x"44";
             when "00001001011010" => D <= x"45";
             when "00001001011011" => D <= x"46";
             when "00001001011100" => D <= x"47";
             when "00001001011101" => D <= x"48";
             when "00001001011110" => D <= x"49";
             when "00001001011111" => D <= x"4A";
             when "00001001100000" => D <= x"4B";
             when "00001001100001" => D <= x"4C";
             when "00001001100010" => D <= x"4D";
             when "00001001100011" => D <= x"4E";
             when "00001001100100" => D <= x"4F";
             when "00001001100101" => D <= x"50";
             when "00001001100110" => D <= x"51";
             when "00001001100111" => D <= x"52";
             when "00001001101000" => D <= x"53";
             when "00001001101001" => D <= x"54";
             when "00001001101010" => D <= x"55";
             when "00001001101011" => D <= x"56";
             when "00001001101100" => D <= x"57";
             when "00001001101101" => D <= x"58";
             when "00001001101110" => D <= x"59";
             when "00001001101111" => D <= x"5A";
             when "00001001110000" => D <= x"00";
             when "00001001110001" => D <= x"20";
             when "00001001110010" => D <= x"20";
             when "00001001110011" => D <= x"61";
             when "00001001110100" => D <= x"62";
             when "00001001110101" => D <= x"63";
             when "00001001110110" => D <= x"64";
             when "00001001110111" => D <= x"65";
             when "00001001111000" => D <= x"66";
             when "00001001111001" => D <= x"67";
             when "00001001111010" => D <= x"68";
             when "00001001111011" => D <= x"69";
             when "00001001111100" => D <= x"6A";
             when "00001001111101" => D <= x"6B";
             when "00001001111110" => D <= x"6C";
             when "00001001111111" => D <= x"6D";
             when "00001010000000" => D <= x"6E";
             when "00001010000001" => D <= x"6F";
             when "00001010000010" => D <= x"70";
             when "00001010000011" => D <= x"71";
             when "00001010000100" => D <= x"72";
             when "00001010000101" => D <= x"73";
             when "00001010000110" => D <= x"74";
             when "00001010000111" => D <= x"75";
             when "00001010001000" => D <= x"76";
             when "00001010001001" => D <= x"77";
             when "00001010001010" => D <= x"78";
             when "00001010001011" => D <= x"79";
             when "00001010001100" => D <= x"7A";
             when "00001010001101" => D <= x"00";
             when "00001010001110" => D <= x"20";
             when "00001010001111" => D <= x"20";
             when "00001010010000" => D <= x"20";
             when "00001010010001" => D <= x"20";
             when "00001010010010" => D <= x"20";
             when "00001010010011" => D <= x"20";
             when "00001010010100" => D <= x"20";
             when "00001010010101" => D <= x"20";
             when "00001010010110" => D <= x"20";
             when "00001010010111" => D <= x"30";
             when "00001010011000" => D <= x"31";
             when "00001010011001" => D <= x"32";
             when "00001010011010" => D <= x"33";
             when "00001010011011" => D <= x"34";
             when "00001010011100" => D <= x"35";
             when "00001010011101" => D <= x"36";
             when "00001010011110" => D <= x"37";
             when "00001010011111" => D <= x"38";
             when "00001010100000" => D <= x"39";
             when "00001010100001" => D <= x"00";
             when "00001010100010" => D <= x"02";
             when "00001010100011" => D <= x"03";
             when "00001010100100" => D <= x"04";
             when "00001010100101" => D <= x"0B";
             when "00001010100110" => D <= x"0C";
             when "00001010100111" => D <= x"0D";
             when "00001010101000" => D <= x"0E";
             when "00001010101001" => D <= x"12";
             when "00001010101010" => D <= x"18";
             when "00001010101011" => D <= x"19";
             when "00001010101100" => D <= x"1A";
             when "00001010101101" => D <= x"1B";
             when "00001010101110" => D <= x"E8";
             when "00001010101111" => D <= x"E9";
             when "00001010110000" => D <= x"EB";
             when "00001010110001" => D <= x"BB";
             when "00001010110010" => D <= x"BC";
             when "00001010110011" => D <= x"8A";
             when "00001010110100" => D <= x"86";
             when "00001010110101" => D <= x"87";
             when "00001010110110" => D <= x"81";
             when "00001010110111" => D <= x"80";
             when "00001010111000" => D <= x"01";
             when "00001010111001" => D <= x"06";
             when "00001010111010" => D <= x"07";
             when "00001010111011" => D <= x"08";
             when "00001010111100" => D <= x"09";
             when "00001010111101" => D <= x"0A";
             when "00001010111110" => D <= x"1D";
             when "00001010111111" => D <= x"1F";
             when "00001011000000" => D <= x"00";
             when "00001011000001" => D <= x"C9";
             when "00001011000010" => D <= x"CD";
             when "00001011000011" => D <= x"CD";
             when "00001011000100" => D <= x"CD";
             when "00001011000101" => D <= x"CD";
             when "00001011000110" => D <= x"CD";
             when "00001011000111" => D <= x"CD";
             when "00001011001000" => D <= x"CD";
             when "00001011001001" => D <= x"CD";
             when "00001011001010" => D <= x"CD";
             when "00001011001011" => D <= x"CD";
             when "00001011001100" => D <= x"CD";
             when "00001011001101" => D <= x"CD";
             when "00001011001110" => D <= x"CD";
             when "00001011001111" => D <= x"CD";
             when "00001011010000" => D <= x"CD";
             when "00001011010001" => D <= x"CD";
             when "00001011010010" => D <= x"CD";
             when "00001011010011" => D <= x"CD";
             when "00001011010100" => D <= x"CD";
             when "00001011010101" => D <= x"CD";
             when "00001011010110" => D <= x"CD";
             when "00001011010111" => D <= x"CD";
             when "00001011011000" => D <= x"CD";
             when "00001011011001" => D <= x"CD";
             when "00001011011010" => D <= x"CD";
             when "00001011011011" => D <= x"CD";
             when "00001011011100" => D <= x"CD";
             when "00001011011101" => D <= x"CD";
             when "00001011011110" => D <= x"CD";
             when "00001011011111" => D <= x"CD";
             when "00001011100000" => D <= x"BB";
             when "00001011100001" => D <= x"00";
             when "00001011100010" => D <= x"C8";
             when "00001011100011" => D <= x"CD";
             when "00001011100100" => D <= x"CD";
             when "00001011100101" => D <= x"CD";
             when "00001011100110" => D <= x"CD";
             when "00001011100111" => D <= x"CD";
             when "00001011101000" => D <= x"CD";
             when "00001011101001" => D <= x"CD";
             when "00001011101010" => D <= x"CD";
             when "00001011101011" => D <= x"CD";
             when "00001011101100" => D <= x"CD";
             when "00001011101101" => D <= x"CD";
             when "00001011101110" => D <= x"CD";
             when "00001011101111" => D <= x"CD";
             when "00001011110000" => D <= x"CD";
             when "00001011110001" => D <= x"CD";
             when "00001011110010" => D <= x"CD";
             when "00001011110011" => D <= x"CD";
             when "00001011110100" => D <= x"CD";
             when "00001011110101" => D <= x"CD";
             when "00001011110110" => D <= x"CD";
             when "00001011110111" => D <= x"CD";
             when "00001011111000" => D <= x"CD";
             when "00001011111001" => D <= x"CD";
             when "00001011111010" => D <= x"CD";
             when "00001011111011" => D <= x"CD";
             when "00001011111100" => D <= x"CD";
             when "00001011111101" => D <= x"CD";
             when "00001011111110" => D <= x"CD";
             when "00001011111111" => D <= x"CD";
             when "00001100000000" => D <= x"CD";
             when "00001100000001" => D <= x"BC";
             when "00001100000010" => D <= x"00";
             when "00001100000011" => D <= x"BA";
             when "00001100000100" => D <= x"20";
             when "00001100000101" => D <= x"20";
             when "00001100000110" => D <= x"20";
             when "00001100000111" => D <= x"20";
             when "00001100001000" => D <= x"20";
             when "00001100001001" => D <= x"20";
             when "00001100001010" => D <= x"20";
             when "00001100001011" => D <= x"20";
             when "00001100001100" => D <= x"20";
             when "00001100001101" => D <= x"20";
             when "00001100001110" => D <= x"20";
             when "00001100001111" => D <= x"20";
             when "00001100010000" => D <= x"20";
             when "00001100010001" => D <= x"20";
             when "00001100010010" => D <= x"20";
             when "00001100010011" => D <= x"20";
             when "00001100010100" => D <= x"20";
             when "00001100010101" => D <= x"20";
             when "00001100010110" => D <= x"20";
             when "00001100010111" => D <= x"20";
             when "00001100011000" => D <= x"20";
             when "00001100011001" => D <= x"20";
             when "00001100011010" => D <= x"20";
             when "00001100011011" => D <= x"20";
             when "00001100011100" => D <= x"20";
             when "00001100011101" => D <= x"20";
             when "00001100011110" => D <= x"20";
             when "00001100011111" => D <= x"20";
             when "00001100100000" => D <= x"20";
             when "00001100100001" => D <= x"20";
             when "00001100100010" => D <= x"BA";
             when "00001100100011" => D <= x"00";
             when "00001100100100" => D <= x"20";
             when "00001100100101" => D <= x"20";
             when "00001100100110" => D <= x"20";
             when "00001100100111" => D <= x"5A";
             when "00001100101000" => D <= x"38";
             when "00001100101001" => D <= x"30";
             when "00001100101010" => D <= x"20";
             when "00001100101011" => D <= x"53";
             when "00001100101100" => D <= x"59";
             when "00001100101101" => D <= x"53";
             when "00001100101110" => D <= x"54";
             when "00001100101111" => D <= x"45";
             when "00001100110000" => D <= x"4D";
             when "00001100110001" => D <= x"20";
             when "00001100110010" => D <= x"20";
             when "00001100110011" => D <= x"20";
             when "00001100110100" => D <= x"20";
             when "00001100110101" => D <= x"52";
             when "00001100110110" => D <= x"4F";
             when "00001100110111" => D <= x"4E";
             when "00001100111000" => D <= x"49";
             when "00001100111001" => D <= x"56";
             when "00001100111010" => D <= x"4F";
             when "00001100111011" => D <= x"4E";
             when "00001100111100" => D <= x"20";
             when "00001100111101" => D <= x"20";
             when "00001100111110" => D <= x"43";
             when "00001100111111" => D <= x"4F";
             when "00001101000000" => D <= x"53";
             when "00001101000001" => D <= x"54";
             when "00001101000010" => D <= x"41";
             when "00001101000011" => D <= x"20";
             when "00001101000100" => D <= x"00";
             when "00001101000101" => D <= x"44";
             when "00001101000110" => D <= x"45";
             when "00001101000111" => D <= x"31";
             when "00001101001000" => D <= x"20";
             when "00001101001001" => D <= x"56";
             when "00001101001010" => D <= x"65";
             when "00001101001011" => D <= x"72";
             when "00001101001100" => D <= x"73";
             when "00001101001101" => D <= x"69";
             when "00001101001110" => D <= x"6F";
             when "00001101001111" => D <= x"6E";
             when "00001101010000" => D <= x"00";
             when "00001101010001" => D <= x"53";
             when "00001101010010" => D <= x"33";
             when "00001101010011" => D <= x"45";
             when "00001101010100" => D <= x"20";
             when "00001101010101" => D <= x"56";
             when "00001101010110" => D <= x"65";
             when "00001101010111" => D <= x"72";
             when "00001101011000" => D <= x"73";
             when "00001101011001" => D <= x"69";
             when "00001101011010" => D <= x"6F";
             when "00001101011011" => D <= x"6E";
             when "00001101011100" => D <= x"00";
             when others => D <= "ZZZZZZZZ";
        end case;
 end if;
end process;
end;
