library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
	port(
		Clk		: in std_logic;
		A		: in std_logic_vector(15 downto 0);
		D		: out std_logic_vector(7 downto 0)
	);
end rom;

architecture rtl of rom is
begin

process (Clk)
begin
 if Clk'event and Clk = '1' then
	case A is
             when x"0000" => D <= x"31";
             when x"0001" => D <= x"FF";
             when x"0002" => D <= x"FF";
             when x"0003" => D <= x"11";
             when x"0004" => D <= x"33";
             when x"0005" => D <= x"20";
             when x"0006" => D <= x"21";
             when x"0007" => D <= x"B7";
             when x"0008" => D <= x"00";
             when x"0009" => D <= x"CD";
             when x"000A" => D <= x"A6";
             when x"000B" => D <= x"00";
             when x"000C" => D <= x"11";
             when x"000D" => D <= x"5B";
             when x"000E" => D <= x"20";
             when x"000F" => D <= x"21";
             when x"0010" => D <= x"CA";
             when x"0011" => D <= x"00";
             when x"0012" => D <= x"CD";
             when x"0013" => D <= x"A6";
             when x"0014" => D <= x"00";
             when x"0015" => D <= x"DB";
             when x"0016" => D <= x"20";
             when x"0017" => D <= x"32";
             when x"0018" => D <= x"00";
             when x"0019" => D <= x"E0";
             when x"001A" => D <= x"CD";
             when x"001B" => D <= x"96";
             when x"001C" => D <= x"00";
             when x"001D" => D <= x"11";
             when x"001E" => D <= x"00";
             when x"001F" => D <= x"20";
             when x"0020" => D <= x"01";
             when x"0021" => D <= x"B0";
             when x"0022" => D <= x"04";
             when x"0023" => D <= x"CD";
             when x"0024" => D <= x"AE";
             when x"0025" => D <= x"00";
             when x"0026" => D <= x"FE";
             when x"0027" => D <= x"41";
             when x"0028" => D <= x"28";
             when x"0029" => D <= x"0B";
             when x"002A" => D <= x"D3";
             when x"002B" => D <= x"11";
             when x"002C" => D <= x"12";
             when x"002D" => D <= x"13";
             when x"002E" => D <= x"0B";
             when x"002F" => D <= x"78";
             when x"0030" => D <= x"B1";
             when x"0031" => D <= x"28";
             when x"0032" => D <= x"EA";
             when x"0033" => D <= x"18";
             when x"0034" => D <= x"EE";
             when x"0035" => D <= x"21";
             when x"0036" => D <= x"00";
             when x"0037" => D <= x"40";
             when x"0038" => D <= x"3E";
             when x"0039" => D <= x"00";
             when x"003A" => D <= x"77";
             when x"003B" => D <= x"23";
             when x"003C" => D <= x"3C";
             when x"003D" => D <= x"20";
             when x"003E" => D <= x"FB";
             when x"003F" => D <= x"3E";
             when x"0040" => D <= x"01";
             when x"0041" => D <= x"D3";
             when x"0042" => D <= x"01";
             when x"0043" => D <= x"CD";
             when x"0044" => D <= x"88";
             when x"0045" => D <= x"00";
             when x"0046" => D <= x"CD";
             when x"0047" => D <= x"88";
             when x"0048" => D <= x"00";
             when x"0049" => D <= x"CD";
             when x"004A" => D <= x"88";
             when x"004B" => D <= x"00";
             when x"004C" => D <= x"CD";
             when x"004D" => D <= x"75";
             when x"004E" => D <= x"00";
             when x"004F" => D <= x"CD";
             when x"0050" => D <= x"88";
             when x"0051" => D <= x"00";
             when x"0052" => D <= x"CD";
             when x"0053" => D <= x"75";
             when x"0054" => D <= x"00";
             when x"0055" => D <= x"21";
             when x"0056" => D <= x"00";
             when x"0057" => D <= x"40";
             when x"0058" => D <= x"7C";
             when x"0059" => D <= x"D3";
             when x"005A" => D <= x"11";
             when x"005B" => D <= x"7D";
             when x"005C" => D <= x"D3";
             when x"005D" => D <= x"10";
             when x"005E" => D <= x"7E";
             when x"005F" => D <= x"D3";
             when x"0060" => D <= x"01";
             when x"0061" => D <= x"CD";
             when x"0062" => D <= x"88";
             when x"0063" => D <= x"00";
             when x"0064" => D <= x"23";
             when x"0065" => D <= x"7E";
             when x"0066" => D <= x"FE";
             when x"0067" => D <= x"FF";
             when x"0068" => D <= x"20";
             when x"0069" => D <= x"EE";
             when x"006A" => D <= x"3E";
             when x"006B" => D <= x"00";
             when x"006C" => D <= x"D3";
             when x"006D" => D <= x"01";
             when x"006E" => D <= x"D3";
             when x"006F" => D <= x"02";
             when x"0070" => D <= x"CD";
             when x"0071" => D <= x"75";
             when x"0072" => D <= x"00";
             when x"0073" => D <= x"18";
             when x"0074" => D <= x"A5";
             when x"0075" => D <= x"CD";
             when x"0076" => D <= x"88";
             when x"0077" => D <= x"00";
             when x"0078" => D <= x"DB";
             when x"0079" => D <= x"30";
             when x"007A" => D <= x"D3";
             when x"007B" => D <= x"10";
             when x"007C" => D <= x"FE";
             when x"007D" => D <= x"0E";
             when x"007E" => D <= x"20";
             when x"007F" => D <= x"F5";
             when x"0080" => D <= x"C9";
             when x"0081" => D <= x"3A";
             when x"0082" => D <= x"00";
             when x"0083" => D <= x"E0";
             when x"0084" => D <= x"3D";
             when x"0085" => D <= x"20";
             when x"0086" => D <= x"FD";
             when x"0087" => D <= x"C9";
             when x"0088" => D <= x"3A";
             when x"0089" => D <= x"00";
             when x"008A" => D <= x"E0";
             when x"008B" => D <= x"F5";
             when x"008C" => D <= x"3E";
             when x"008D" => D <= x"FF";
             when x"008E" => D <= x"3D";
             when x"008F" => D <= x"20";
             when x"0090" => D <= x"FD";
             when x"0091" => D <= x"F1";
             when x"0092" => D <= x"3D";
             when x"0093" => D <= x"20";
             when x"0094" => D <= x"F6";
             when x"0095" => D <= x"C9";
             when x"0096" => D <= x"21";
             when x"0097" => D <= x"00";
             when x"0098" => D <= x"20";
             when x"0099" => D <= x"11";
             when x"009A" => D <= x"B0";
             when x"009B" => D <= x"04";
             when x"009C" => D <= x"3E";
             when x"009D" => D <= x"20";
             when x"009E" => D <= x"77";
             when x"009F" => D <= x"23";
             when x"00A0" => D <= x"1B";
             when x"00A1" => D <= x"7A";
             when x"00A2" => D <= x"B3";
             when x"00A3" => D <= x"20";
             when x"00A4" => D <= x"F7";
             when x"00A5" => D <= x"C9";
             when x"00A6" => D <= x"7E";
             when x"00A7" => D <= x"B7";
             when x"00A8" => D <= x"C8";
             when x"00A9" => D <= x"12";
             when x"00AA" => D <= x"23";
             when x"00AB" => D <= x"13";
             when x"00AC" => D <= x"18";
             when x"00AD" => D <= x"F8";
             when x"00AE" => D <= x"CD";
             when x"00AF" => D <= x"88";
             when x"00B0" => D <= x"00";
             when x"00B1" => D <= x"DB";
             when x"00B2" => D <= x"80";
             when x"00B3" => D <= x"B7";
             when x"00B4" => D <= x"28";
             when x"00B5" => D <= x"F8";
             when x"00B6" => D <= x"C9";
             when x"00B7" => D <= x"5A";
             when x"00B8" => D <= x"38";
             when x"00B9" => D <= x"30";
             when x"00BA" => D <= x"20";
             when x"00BB" => D <= x"53";
             when x"00BC" => D <= x"59";
             when x"00BD" => D <= x"53";
             when x"00BE" => D <= x"54";
             when x"00BF" => D <= x"45";
             when x"00C0" => D <= x"4D";
             when x"00C1" => D <= x"20";
             when x"00C2" => D <= x"4F";
             when x"00C3" => D <= x"4E";
             when x"00C4" => D <= x"20";
             when x"00C5" => D <= x"43";
             when x"00C6" => D <= x"48";
             when x"00C7" => D <= x"49";
             when x"00C8" => D <= x"50";
             when x"00C9" => D <= x"00";
             when x"00CA" => D <= x"52";
             when x"00CB" => D <= x"4F";
             when x"00CC" => D <= x"4E";
             when x"00CD" => D <= x"49";
             when x"00CE" => D <= x"56";
             when x"00CF" => D <= x"4F";
             when x"00D0" => D <= x"4E";
             when x"00D1" => D <= x"20";
             when x"00D2" => D <= x"43";
             when x"00D3" => D <= x"4F";
             when x"00D4" => D <= x"53";
             when x"00D5" => D <= x"54";
             when x"00D6" => D <= x"41";
             when x"00D7" => D <= x"20";
             when x"00D8" => D <= x"32";
             when x"00D9" => D <= x"30";
             when x"00DA" => D <= x"30";
             when x"00DB" => D <= x"38";
             when x"00DC" => D <= x"00";
             when others => D <= x"00";
	end case;
 end if;
end process;
end;
